MOSFET Half Bridge Driver

.INCLUDE BC847.prm
.INCLUDE BC857.prm
.INCLUDE IRF7303.prm
.INCLUDE IRF7304.prm

R1 1   2  100K
R2 100 3   22K
R3 100 6   22K
R4   5 6    1K



*    C B E
Q1   3 1 5 QBC847
Q2   6 2 0 QBC847
Q3 100 3 4 QBC847

.model D1N4148  D(IS=35p RS=64m N=1.24 TT=5n CJO=4p M=0.285 VJ=0.6 BV=75)
.model ZDIODE15 D(BV=15V IBV=17m )
D2   4 3 D1N4148
D3   0 6 ZDIODE15

* M4   10 4 100 100
* M5   11 6   0   0
X4   10 4 100 irf7304 
X5   11 6   0 auirf7303q

VSUPPLY   100  0 12V
VDUMMY    10  11  0V
* VCONTROL  1    0  PULSE(0.1 1.7 0 1ns 1ns 1ms 1ms)
VCONTROL  1    0  SIN(0.6VOFF 0.6VPEAK   10HZ)

.END
